library verilog;
use verilog.vl_types.all;
entity test1_tb is
end test1_tb;
