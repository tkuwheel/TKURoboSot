library verilog;
use verilog.vl_types.all;
entity Crc16_tb is
end Crc16_tb;
