library verilog;
use verilog.vl_types.all;
entity Serial2CMD_tb is
end Serial2CMD_tb;
